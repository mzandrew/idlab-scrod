--*********************************************************************************
-- Indiana University
-- Center for Exploration of Energy and Matter (CEEM)
--
-- Project: Belle-II
--
-- Author:  Brandon Kunkler
--
-- Date:    06/05/2014
--
--*********************************************************************************
-- Description:
-- Test bench for time order entity. Uses TDC entity as stimulus. Stimulus can be
-- generated by a counter or a pseudo-random noise generator.
--
-- Deficiencies:
-- Need a more clever way of generating separately for each channel and more slowly.
--*********************************************************************************

library ieee;
    use ieee.std_logic_1164.all;
--    use ieee.math_real.all;
--     use ieee.numeric_std.all;
    use ieee.std_logic_unsigned.all;
    use ieee.std_logic_textio.all;
library work;
    use work.time_order_pkg.all;
    use work.tdc_pkg.all;


entity time_order_tb is
end time_order_tb;

architecture behave of time_order_tb is

    component tdc is
    port(
    -- Inputs -----------------------------
        tdc_clk                     : in std_logic;
        ce                          : in std_logic_vector(1 to 4);
        reset                       : in std_logic;
        tdc_clr                     : in std_logic;
        tb                          : in tb_vec_type;
        tb16                        : in std_logic_vector(1 to TDC_NUM_CHAN);
        fifo_re                     : in std_logic_vector(1 to TDC_NUM_CHAN);
    -- Outputs -----------------------------
        fifo_ept                    : out std_logic_vector(1 to TDC_NUM_CHAN);
        tdc_dout                    : out tdc_dout_type);
    end component;

    component time_order is
        port(
        clk                         : in std_logic;
        ce                          : in std_logic;
        reset                       : in std_logic;
        dst_full                    : in std_logic;
        src_epty                    : in std_logic_vector(1 to TO_NUM_LANES);
        din                         : in tdc_dout_type;
        src_re                      : out std_logic_vector(1 to TO_NUM_LANES);
        dst_we                      : out std_logic;
        dout                        : out std_logic_vector(TO_WIDTH-1 downto 0));
    end component;

    component tdc_stim is
    generic(
        USE_PRNG                    : std_logic);
    port(
        clk                         : in std_logic;
        ce                          : in std_logic;
        stim_enable                 : in std_logic;        
        run_reset                   : in std_logic;
        tb                          : out std_logic_vector(5 downto 1);
        tb16                        : out std_logic);
    end component;

    constant USE_PRNG               : std_logic                             := '0';
    constant CLKPER                 : time                                  := 4 ns;
    constant CLKHLFPER              : time                                  := CLKPER/2;

    signal clk                      : std_logic                             := '1';
    signal ce                       : std_logic_vector(1 to 6)              := (others => '0');
    signal run_reset                : std_logic                             := '1';    
    signal tb                       : tb_vec_type                           := (others => "00000");
    signal tb16                     : std_logic_vector(1 to TDC_NUM_CHAN)   := (others => '0');
    signal fifo_re                  : std_logic_vector(1 to TDC_NUM_CHAN)   := (others => '0');
    signal fifo_ept                 : std_logic_vector(1 to TDC_NUM_CHAN);
    signal tdc_dout                 : tdc_dout_type;       
    signal dst_we                   : std_logic;
    signal dst_full                 : std_logic                             := '0';
    signal ordered                  : std_logic_vector(TO_WIDTH-1 downto 0);
    
    signal ce_bit                   : std_logic                             := '0';        
    signal ce_cnt                   : std_logic_vector(2 downto 0)          := (others => '1');
    signal full_reg                 : std_logic_vector(15 downto 0);    
    signal lordered                 : std_logic_vector(3 downto 0);--lane
    signal cordered                 : std_logic_vector(3 downto 0);--channel
    signal dordered                 : std_logic_vector(TO_DWIDTH-1 downto 0);    
    signal stim_enable              : std_logic                             := '0';
    signal test                     : std_logic;

begin

    ------------------------------------------------------------
    -- Generate stimulus for each lane separately.
    ------------------------------------------------------------    
    STIM_GEN:
    for I in 1 to TO_NUM_LANES generate
    stim_ins : tdc_stim
    generic map(
        USE_PRNG                    => USE_PRNG)
    port map(                       
        clk                         => clk,
        ce                          => ce(6),
        run_reset                   => run_reset,
        stim_enable                 => stim_enable,
        tb                          => tb(I),
        tb16                        => tb16(I));
    end generate;

    ------------------------------------------------------------
    -- Use TDC for stimulus because doing otherwise requires
    -- too much labor.
    ------------------------------------------------------------
    tdc_ins : tdc
    port map(
    -- Inputs -----------------------------
        tdc_clk                     => clk,
        ce                          => ce(1 to 4),
        reset                       => run_reset,
        tdc_clr                     => run_reset,
        tb                          => tb,
        tb16                        => tb16,
        fifo_re                     => fifo_re,
    -- Outputs -----------------------------
        fifo_ept                    => fifo_ept,
        tdc_dout                    => tdc_dout
    );

    ------------------------------------------------------------
    -- UUT: Time order entity
    ------------------------------------------------------------
    UUT : time_order
    port map(
        clk                         => clk,
        ce                          => ce(5),
        reset                       => run_reset,
        dst_full                    => dst_full,
        src_epty                    => fifo_ept,
        din                         => tdc_dout,
        src_re                      => fifo_re,
        dst_we                      => dst_we,
        dout                        => ordered
    );

    -- Generate clock
    clk <= (not clk) after CLKHLFPER;
    -- Simulate power on reset
    run_reset <= '0' after CLKPER*8;    
    stim_enable <= not run_reset'delayed(CLKPER*12);
    ce <= (others => ce_bit);

    dst_full <= full_reg(5);

    lordered <= ordered(ordered'length-1 downto ordered'length-4);--lane
    cordered <= ordered(ordered'length-5 downto ordered'length-TO_CWIDTH);--channel
    dordered <= ordered(TO_DWIDTH-1 downto 0);--TDC

    --------------------------------------------------------------------------
    -- Generate a psuedo-random shift register for creating a full signal at
    -- different intervals. Provide stimulus that fully verifies time order
    -- circuit by toggling the receiving entities full flag.
    --------------------------------------------------------------------------
    full_pcs : process(run_reset,clk)
    begin
        if run_reset = '1' then
            full_reg <= "0110110010101001";
        else
            if rising_edge(clk) then
                full_reg <= full_reg(14 downto 0) & (full_reg(15) xor full_reg(12));
            end if;
        end if;
    end process;

    --------------------------------------------------------------------------
    -- Generate clock enable.
    --------------------------------------------------------------------------
    ce_cnt_pcs : process(run_reset,clk)
    begin
        if run_reset = '1' then
            ce_cnt <= (others => '0');
        else
            if rising_edge(clk) then
                ce_cnt <= ce_cnt + 1;
            end if;
        end if;
    end process;

    ce2x_pcs : process
    begin
        wait until rising_edge(ce_cnt(0));
            ce_bit <= '1';
        wait for CLKPER;
            ce_bit <= '0';
    end process;

end behave;