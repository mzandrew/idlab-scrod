`timescale 1ns/1ps

/****************************************************************************
	University of Hawaii at Manoa
	Instrumentation Development Lab / GARY S. VARNER
	Watanabe Hall Room 214
	2505 Correa Road
	Honolulu, HI 96822
	Lab: (808) 956-2920
	Fax: (808) 956-2930
	E-mail: idlab@phys.hawaii.edu
	
AND
	
	Pacific Northwest National Laboratory
	902 Battelle Blvd., MS J4-60
	Richland, WA  99352
	
 ****************************************************************************

	Design by:	Lynn Wood, PNNL (lynn.wood@pnnl.gov)
	Started:		11 Jul 2011
	Project:		Belle II iTOP firmware
	
	Description:
		Provides a fixed time delay by using the carry chain of a single 
		column in the FPGA.  To ensure a consistent delay value, the locations
		of each element are constrained to an exact X,Y location in the FPGA.

 ****************************************************************************/


// carry chain automatically generated by gen_carrychain.exe
module SMPL_CARRY_CHAIN(cin, cout);
	input		cin;
	output	cout;
	
	wire	[159:0]	dly;
	
//	assign cout = dly[159];
	assign cout = dly[155];
//	assign cout = dly[151];
//	assign cout = dly[143];
//	assign cout = dly[134];
//	assign cout = dly[127];
//	assign cout = dly[111];
//	assign cout = dly[95];
//	assign cout = dly[79];
//	assign cout = dly[63];


   (* LOC="SLICE_X2Y16" *)  MUXCY_L muxcy00(.LO(dly[ 0]), .CI(    cin), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y17" *)  MUXCY_L muxcy01(.LO(dly[ 1]), .CI(dly[ 0]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y18" *)  MUXCY_L muxcy02(.LO(dly[ 2]), .CI(dly[ 1]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y19" *)  MUXCY_L muxcy03(.LO(dly[ 3]), .CI(dly[ 2]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y20" *)  MUXCY_L muxcy04(.LO(dly[ 4]), .CI(dly[ 3]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y21" *)  MUXCY_L muxcy05(.LO(dly[ 5]), .CI(dly[ 4]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y22" *)  MUXCY_L muxcy06(.LO(dly[ 6]), .CI(dly[ 5]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y23" *)  MUXCY_L muxcy07(.LO(dly[ 7]), .CI(dly[ 6]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y24" *)  MUXCY_L muxcy08(.LO(dly[ 8]), .CI(dly[ 7]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y25" *)  MUXCY_L muxcy09(.LO(dly[ 9]), .CI(dly[ 8]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y26" *)  MUXCY_L muxcy10(.LO(dly[10]), .CI(dly[ 9]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y27" *)  MUXCY_L muxcy11(.LO(dly[11]), .CI(dly[10]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y28" *)  MUXCY_L muxcy12(.LO(dly[12]), .CI(dly[11]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y29" *)  MUXCY_L muxcy13(.LO(dly[13]), .CI(dly[12]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y30" *)  MUXCY_L muxcy14(.LO(dly[14]), .CI(dly[13]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y31" *)  MUXCY_L muxcy15(.LO(dly[15]), .CI(dly[14]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y32" *)  MUXCY_L muxcy16(.LO(dly[16]), .CI(dly[15]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y33" *)  MUXCY_L muxcy17(.LO(dly[17]), .CI(dly[16]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y34" *)  MUXCY_L muxcy18(.LO(dly[18]), .CI(dly[17]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y35" *)  MUXCY_L muxcy19(.LO(dly[19]), .CI(dly[18]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y36" *)  MUXCY_L muxcy20(.LO(dly[20]), .CI(dly[19]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y37" *)  MUXCY_L muxcy21(.LO(dly[21]), .CI(dly[20]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y38" *)  MUXCY_L muxcy22(.LO(dly[22]), .CI(dly[21]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y39" *)  MUXCY_L muxcy23(.LO(dly[23]), .CI(dly[22]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y40" *)  MUXCY_L muxcy24(.LO(dly[24]), .CI(dly[23]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y41" *)  MUXCY_L muxcy25(.LO(dly[25]), .CI(dly[24]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y42" *)  MUXCY_L muxcy26(.LO(dly[26]), .CI(dly[25]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y43" *)  MUXCY_L muxcy27(.LO(dly[27]), .CI(dly[26]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y44" *)  MUXCY_L muxcy28(.LO(dly[28]), .CI(dly[27]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y45" *)  MUXCY_L muxcy29(.LO(dly[29]), .CI(dly[28]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y46" *)  MUXCY_L muxcy30(.LO(dly[30]), .CI(dly[29]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y47" *)  MUXCY_L muxcy31(.LO(dly[31]), .CI(dly[30]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y48" *)  MUXCY_L muxcy32(.LO(dly[32]), .CI(dly[31]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y49" *)  MUXCY_L muxcy33(.LO(dly[33]), .CI(dly[32]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y50" *)  MUXCY_L muxcy34(.LO(dly[34]), .CI(dly[33]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y51" *)  MUXCY_L muxcy35(.LO(dly[35]), .CI(dly[34]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y52" *)  MUXCY_L muxcy36(.LO(dly[36]), .CI(dly[35]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y53" *)  MUXCY_L muxcy37(.LO(dly[37]), .CI(dly[36]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y54" *)  MUXCY_L muxcy38(.LO(dly[38]), .CI(dly[37]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y55" *)  MUXCY_L muxcy39(.LO(dly[39]), .CI(dly[38]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y56" *)  MUXCY_L muxcy40(.LO(dly[40]), .CI(dly[39]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y57" *)  MUXCY_L muxcy41(.LO(dly[41]), .CI(dly[40]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y58" *)  MUXCY_L muxcy42(.LO(dly[42]), .CI(dly[41]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y59" *)  MUXCY_L muxcy43(.LO(dly[43]), .CI(dly[42]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y60" *)  MUXCY_L muxcy44(.LO(dly[44]), .CI(dly[43]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y61" *)  MUXCY_L muxcy45(.LO(dly[45]), .CI(dly[44]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y62" *)  MUXCY_L muxcy46(.LO(dly[46]), .CI(dly[45]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y63" *)  MUXCY_L muxcy47(.LO(dly[47]), .CI(dly[46]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y64" *)  MUXCY_L muxcy48(.LO(dly[48]), .CI(dly[47]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y65" *)  MUXCY_L muxcy49(.LO(dly[49]), .CI(dly[48]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y66" *)  MUXCY_L muxcy50(.LO(dly[50]), .CI(dly[49]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y67" *)  MUXCY_L muxcy51(.LO(dly[51]), .CI(dly[50]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y68" *)  MUXCY_L muxcy52(.LO(dly[52]), .CI(dly[51]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y69" *)  MUXCY_L muxcy53(.LO(dly[53]), .CI(dly[52]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y70" *)  MUXCY_L muxcy54(.LO(dly[54]), .CI(dly[53]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y71" *)  MUXCY_L muxcy55(.LO(dly[55]), .CI(dly[54]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y72" *)  MUXCY_L muxcy56(.LO(dly[56]), .CI(dly[55]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y73" *)  MUXCY_L muxcy57(.LO(dly[57]), .CI(dly[56]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y74" *)  MUXCY_L muxcy58(.LO(dly[58]), .CI(dly[57]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y75" *)  MUXCY_L muxcy59(.LO(dly[59]), .CI(dly[58]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y76" *)  MUXCY_L muxcy60(.LO(dly[60]), .CI(dly[59]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y77" *)  MUXCY_L muxcy61(.LO(dly[61]), .CI(dly[60]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y78" *)  MUXCY_L muxcy62(.LO(dly[62]), .CI(dly[61]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y79" *)  MUXCY_L muxcy63(.LO(dly[63]), .CI(dly[62]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y80" *)  MUXCY_L muxcy64(.LO(dly[64]), .CI(dly[63]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y81" *)  MUXCY_L muxcy65(.LO(dly[65]), .CI(dly[64]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y82" *)  MUXCY_L muxcy66(.LO(dly[66]), .CI(dly[65]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y83" *)  MUXCY_L muxcy67(.LO(dly[67]), .CI(dly[66]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y84" *)  MUXCY_L muxcy68(.LO(dly[68]), .CI(dly[67]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y85" *)  MUXCY_L muxcy69(.LO(dly[69]), .CI(dly[68]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y86" *)  MUXCY_L muxcy70(.LO(dly[70]), .CI(dly[69]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y87" *)  MUXCY_L muxcy71(.LO(dly[71]), .CI(dly[70]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y88" *)  MUXCY_L muxcy72(.LO(dly[72]), .CI(dly[71]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y89" *)  MUXCY_L muxcy73(.LO(dly[73]), .CI(dly[72]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y90" *)  MUXCY_L muxcy74(.LO(dly[74]), .CI(dly[73]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y91" *)  MUXCY_L muxcy75(.LO(dly[75]), .CI(dly[74]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y92" *)  MUXCY_L muxcy76(.LO(dly[76]), .CI(dly[75]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y93" *)  MUXCY_L muxcy77(.LO(dly[77]), .CI(dly[76]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y94" *)  MUXCY_L muxcy78(.LO(dly[78]), .CI(dly[77]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y95" *)  MUXCY_L muxcy79(.LO(dly[79]), .CI(dly[78]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y96" *)  MUXCY_L muxcy80(.LO(dly[80]), .CI(dly[79]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y97" *)  MUXCY_L muxcy81(.LO(dly[81]), .CI(dly[80]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y98" *)  MUXCY_L muxcy82(.LO(dly[82]), .CI(dly[81]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y99" *)  MUXCY_L muxcy83(.LO(dly[83]), .CI(dly[82]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y100" *)  MUXCY_L muxcy84(.LO(dly[84]), .CI(dly[83]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y101" *)  MUXCY_L muxcy85(.LO(dly[85]), .CI(dly[84]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y102" *)  MUXCY_L muxcy86(.LO(dly[86]), .CI(dly[85]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y103" *)  MUXCY_L muxcy87(.LO(dly[87]), .CI(dly[86]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y104" *)  MUXCY_L muxcy88(.LO(dly[88]), .CI(dly[87]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y105" *)  MUXCY_L muxcy89(.LO(dly[89]), .CI(dly[88]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y106" *)  MUXCY_L muxcy90(.LO(dly[90]), .CI(dly[89]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y107" *)  MUXCY_L muxcy91(.LO(dly[91]), .CI(dly[90]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y108" *)  MUXCY_L muxcy92(.LO(dly[92]), .CI(dly[91]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y109" *)  MUXCY_L muxcy93(.LO(dly[93]), .CI(dly[92]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y110" *)  MUXCY_L muxcy94(.LO(dly[94]), .CI(dly[93]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y111" *)  MUXCY_L muxcy95(.LO(dly[95]), .CI(dly[94]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y112" *)  MUXCY_L muxcy96(.LO(dly[96]), .CI(dly[95]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y113" *)  MUXCY_L muxcy97(.LO(dly[97]), .CI(dly[96]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y114" *)  MUXCY_L muxcy98(.LO(dly[98]), .CI(dly[97]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y115" *)  MUXCY_L muxcy99(.LO(dly[99]), .CI(dly[98]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y116" *)  MUXCY_L muxcy100(.LO(dly[100]), .CI(dly[99]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y117" *)  MUXCY_L muxcy101(.LO(dly[101]), .CI(dly[100]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y118" *)  MUXCY_L muxcy102(.LO(dly[102]), .CI(dly[101]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y119" *)  MUXCY_L muxcy103(.LO(dly[103]), .CI(dly[102]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y120" *)  MUXCY_L muxcy104(.LO(dly[104]), .CI(dly[103]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y121" *)  MUXCY_L muxcy105(.LO(dly[105]), .CI(dly[104]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y122" *)  MUXCY_L muxcy106(.LO(dly[106]), .CI(dly[105]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y123" *)  MUXCY_L muxcy107(.LO(dly[107]), .CI(dly[106]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y124" *)  MUXCY_L muxcy108(.LO(dly[108]), .CI(dly[107]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y125" *)  MUXCY_L muxcy109(.LO(dly[109]), .CI(dly[108]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y126" *)  MUXCY_L muxcy110(.LO(dly[110]), .CI(dly[109]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y127" *)  MUXCY_L muxcy111(.LO(dly[111]), .CI(dly[110]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y128" *)  MUXCY_L muxcy112(.LO(dly[112]), .CI(dly[111]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y129" *)  MUXCY_L muxcy113(.LO(dly[113]), .CI(dly[112]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y130" *)  MUXCY_L muxcy114(.LO(dly[114]), .CI(dly[113]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y131" *)  MUXCY_L muxcy115(.LO(dly[115]), .CI(dly[114]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y132" *)  MUXCY_L muxcy116(.LO(dly[116]), .CI(dly[115]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y133" *)  MUXCY_L muxcy117(.LO(dly[117]), .CI(dly[116]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y134" *)  MUXCY_L muxcy118(.LO(dly[118]), .CI(dly[117]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y135" *)  MUXCY_L muxcy119(.LO(dly[119]), .CI(dly[118]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y136" *)  MUXCY_L muxcy120(.LO(dly[120]), .CI(dly[119]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y137" *)  MUXCY_L muxcy121(.LO(dly[121]), .CI(dly[120]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y138" *)  MUXCY_L muxcy122(.LO(dly[122]), .CI(dly[121]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y139" *)  MUXCY_L muxcy123(.LO(dly[123]), .CI(dly[122]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y140" *)  MUXCY_L muxcy124(.LO(dly[124]), .CI(dly[123]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y141" *)  MUXCY_L muxcy125(.LO(dly[125]), .CI(dly[124]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y142" *)  MUXCY_L muxcy126(.LO(dly[126]), .CI(dly[125]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y143" *)  MUXCY_L muxcy127(.LO(dly[127]), .CI(dly[126]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y144" *)  MUXCY_L muxcy128(.LO(dly[128]), .CI(dly[127]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y145" *)  MUXCY_L muxcy129(.LO(dly[129]), .CI(dly[128]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y146" *)  MUXCY_L muxcy130(.LO(dly[130]), .CI(dly[129]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y147" *)  MUXCY_L muxcy131(.LO(dly[131]), .CI(dly[130]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y148" *)  MUXCY_L muxcy132(.LO(dly[132]), .CI(dly[131]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y149" *)  MUXCY_L muxcy133(.LO(dly[133]), .CI(dly[132]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y150" *)  MUXCY_L muxcy134(.LO(dly[134]), .CI(dly[133]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y151" *)  MUXCY_L muxcy135(.LO(dly[135]), .CI(dly[134]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y152" *)  MUXCY_L muxcy136(.LO(dly[136]), .CI(dly[135]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y153" *)  MUXCY_L muxcy137(.LO(dly[137]), .CI(dly[136]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y154" *)  MUXCY_L muxcy138(.LO(dly[138]), .CI(dly[137]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y155" *)  MUXCY_L muxcy139(.LO(dly[139]), .CI(dly[138]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y156" *)  MUXCY_L muxcy140(.LO(dly[140]), .CI(dly[139]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y157" *)  MUXCY_L muxcy141(.LO(dly[141]), .CI(dly[140]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y158" *)  MUXCY_L muxcy142(.LO(dly[142]), .CI(dly[141]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y159" *)  MUXCY_L muxcy143(.LO(dly[143]), .CI(dly[142]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y160" *)  MUXCY_L muxcy144(.LO(dly[144]), .CI(dly[143]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y161" *)  MUXCY_L muxcy145(.LO(dly[145]), .CI(dly[144]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y162" *)  MUXCY_L muxcy146(.LO(dly[146]), .CI(dly[145]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y163" *)  MUXCY_L muxcy147(.LO(dly[147]), .CI(dly[146]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y164" *)  MUXCY_L muxcy148(.LO(dly[148]), .CI(dly[147]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y165" *)  MUXCY_L muxcy149(.LO(dly[149]), .CI(dly[148]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y166" *)  MUXCY_L muxcy150(.LO(dly[150]), .CI(dly[149]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y167" *)  MUXCY_L muxcy151(.LO(dly[151]), .CI(dly[150]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y168" *)  MUXCY_L muxcy152(.LO(dly[152]), .CI(dly[151]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y169" *)  MUXCY_L muxcy153(.LO(dly[153]), .CI(dly[152]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y170" *)  MUXCY_L muxcy154(.LO(dly[154]), .CI(dly[153]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y171" *)  MUXCY_L muxcy155(.LO(dly[155]), .CI(dly[154]), .DI(1'b0), .S(1'b1));
/*
   (* LOC="SLICE_X2Y172" *)  MUXCY_L muxcy156(.LO(dly[156]), .CI(dly[155]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y173" *)  MUXCY_L muxcy157(.LO(dly[157]), .CI(dly[156]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y174" *)  MUXCY_L muxcy158(.LO(dly[158]), .CI(dly[157]), .DI(1'b0), .S(1'b1));
   (* LOC="SLICE_X2Y175" *)  MUXCY_L muxcy159(.LO(dly[159]), .CI(dly[158]), .DI(1'b0), .S(1'b1));
*/
endmodule
